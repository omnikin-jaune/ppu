
entity hit_handler is
port (
    i_x        : in vector_pos      (63 downto 0);
    i_y        : in vector_pos      (63 downto 0);
    i_sprite_x : in vector_pos      (63 downto 0);
    i_sprite_y : in vector_pos      (63 downto 0);
    i_en       : in std_logic_vector(63 downto 0);
    i_cc       : in vector_cc       (63 downto 0);

    o_sprite   : out std_logic_vector(5 downto 0);
    o_en       : out std_logic;
) end hit_handler;


architecture behavioral of hit_handler is

    component hit_detector is
    port (
        i_x        : std_logic_vector(8 downto 0);
        i_y        : std_logic_vector(8 downto 0);
        i_sprite_x : std_logic_vector(8 downto 0); 
        i_sprite_y : std_logic_vector(8 downto 0);
        i_en       : std_logic;
        i_cc       : std_logic_vector(5 downto 0);

        o_hit      : std_logic;
    );


    signal s_hits : std_logic_vector(63 downto 0);
    
begin


    -- https://stackoverflow.com/a/13194608
    hit_detector_gen:
    for i in 0 to 63 generate
        hit_detectors: hit_detector
        port map (
            i_x        <= i_x(i),
            i_y        <= i_y(i),
            i_sprite_x <= i_sprite_x(i),
            i_sprite_y <= i_sprite_y(i),
            i_en       <= i_en(i),
            i_cc       <= i_cc(i),
    
            o_hit      <= s_hits(i)
        );
    end generate;


    with s_hits select o_sprite <=
        "00000" when "0000000000000000000000000000000000000000000000000000000000000000",
        "00000" when "0000000000000000000000000000000000000000000000000000000000000001",
        "00000" when "0000000000000000000000000000000000000000000000000000000000000011",
        "00000" when "0000000000000000000000000000000000000000000000000000000000000101",
        "00000" when "0000000000000000000000000000000000000000000000000000000000000111",
        "00000" when "0000000000000000000000000000000000000000000000000000000000001001",
        "00000" when "0000000000000000000000000000000000000000000000000000000000001011",
        "00000" when "0000000000000000000000000000000000000000000000000000000000001101",
        "00000" when "0000000000000000000000000000000000000000000000000000000000001111",
        "00000" when "0000000000000000000000000000000000000000000000000000000000010001",
        "00000" when "0000000000000000000000000000000000000000000000000000000000010011",
        "00000" when "0000000000000000000000000000000000000000000000000000000000010101",
        "00000" when "0000000000000000000000000000000000000000000000000000000000010111",
        "00000" when "0000000000000000000000000000000000000000000000000000000000011001",
        "00000" when "0000000000000000000000000000000000000000000000000000000000011011",
        "00000" when "0000000000000000000000000000000000000000000000000000000000011101",
        "00000" when "0000000000000000000000000000000000000000000000000000000000011111",
        "00000" when "0000000000000000000000000000000000000000000000000000000000100000",
        "00000" when "0000000000000000000000000000000000000000000000000000000000100001",
        "00000" when "0000000000000000000000000000000000000000000000000000000000100010",
        "00000" when "0000000000000000000000000000000000000000000000000000000000100011",
        "00000" when "0000000000000000000000000000000000000000000000000000000000100100",
        "00000" when "0000000000000000000000000000000000000000000000000000000000100101",
        "00000" when "0000000000000000000000000000000000000000000000000000000000100110",
        "00000" when "0000000000000000000000000000000000000000000000000000000000100111",
        "00000" when "0000000000000000000000000000000000000000000000000000000000101000",
        "00000" when "0000000000000000000000000000000000000000000000000000000000101001",
        "00000" when "0000000000000000000000000000000000000000000000000000000000101010",
        "00000" when "0000000000000000000000000000000000000000000000000000000000101011",
        "00000" when "0000000000000000000000000000000000000000000000000000000000101100",
        "00000" when "0000000000000000000000000000000000000000000000000000000000101101",
        "00000" when "0000000000000000000000000000000000000000000000000000000000101110",
        "00000" when "0000000000000000000000000000000000000000000000000000000000101111",
        "00000" when "0000000000000000000000000000000000000000000000000000000000110000",
        "00000" when "0000000000000000000000000000000000000000000000000000000000110001",
        "00000" when "0000000000000000000000000000000000000000000000000000000000110010",
        "00000" when "0000000000000000000000000000000000000000000000000000000000110011",
        "00000" when "0000000000000000000000000000000000000000000000000000000000110100",
        "00000" when "0000000000000000000000000000000000000000000000000000000000110101",
        "00000" when "0000000000000000000000000000000000000000000000000000000000110110",
        "00000" when "0000000000000000000000000000000000000000000000000000000000110111",
        "00000" when "0000000000000000000000000000000000000000000000000000000000111000",
        "00000" when "0000000000000000000000000000000000000000000000000000000000111001",
        "00000" when "0000000000000000000000000000000000000000000000000000000000111010",
        "00000" when "0000000000000000000000000000000000000000000000000000000000111011",
        "00000" when "0000000000000000000000000000000000000000000000000000000000111100",
        "00000" when "0000000000000000000000000000000000000000000000000000000000111101",
        "00000" when "0000000000000000000000000000000000000000000000000000000000111110",
        "00000" when "0000000000000000000000000000000000000000000000000000000000111111",
        "00000" when "0000000000000000000000000000000000000000000000000000000001000000",
        "00000" when "0000000000000000000000000000000000000000000000000000000001000001",
        "00000" when "0000000000000000000000000000000000000000000000000000000001000011",
        "00000" when "0000000000000000000000000000000000000000000000000000000001000101",
        "00000" when "0000000000000000000000000000000000000000000000000000000001000111",
        "00000" when "0000000000000000000000000000000000000000000000000000000001001001",
        "00000" when "0000000000000000000000000000000000000000000000000000000001001011",
        "00000" when "0000000000000000000000000000000000000000000000000000000001001101",
        "00000" when "0000000000000000000000000000000000000000000000000000000001001111",
        "00000" when "0000000000000000000000000000000000000000000000000000000001010001",
        "00000" when "0000000000000000000000000000000000000000000000000000000001010011",
        "00000" when "0000000000000000000000000000000000000000000000000000000001010101",
        "00000" when "0000000000000000000000000000000000000000000000000000000001010111",
        "00000" when "0000000000000000000000000000000000000000000000000000000001011001",
        "00000" when "0000000000000000000000000000000000000000000000000000000001011011",
        "00000" when "0000000000000000000000000000000000000000000000000000000001011101",
        "00000" when "0000000000000000000000000000000000000000000000000000000001011111"
        "00000" when "0000000000000000000000000000000000000000000000000000000001100000",
        "00000" when "0000000000000000000000000000000000000000000000000000000001100001",
        "00000" when "0000000000000000000000000000000000000000000000000000000001100010",
        "00000" when "0000000000000000000000000000000000000000000000000000000001100011",
        "00000" when "0000000000000000000000000000000000000000000000000000000001100100",
        "00000" when "0000000000000000000000000000000000000000000000000000000001100101",
        "00000" when "0000000000000000000000000000000000000000000000000000000001100110",
        "00000" when "0000000000000000000000000000000000000000000000000000000001100111",
        "00000" when "0000000000000000000000000000000000000000000000000000000001101000",
        "00000" when "0000000000000000000000000000000000000000000000000000000001101001",
        "00000" when "0000000000000000000000000000000000000000000000000000000001101010",
        "00000" when "0000000000000000000000000000000000000000000000000000000001101011",
        "00000" when "0000000000000000000000000000000000000000000000000000000001101100",
        "00000" when "0000000000000000000000000000000000000000000000000000000001101101",
        "00000" when "0000000000000000000000000000000000000000000000000000000001101110",
        "00000" when "0000000000000000000000000000000000000000000000000000000001101111",
        "00000" when "0000000000000000000000000000000000000000000000000000000001110000",
        "00000" when "0000000000000000000000000000000000000000000000000000000001110001",
        "00000" when "0000000000000000000000000000000000000000000000000000000001110010",
        "00000" when "0000000000000000000000000000000000000000000000000000000001110011",
        "00000" when "0000000000000000000000000000000000000000000000000000000001110100",
        "00000" when "0000000000000000000000000000000000000000000000000000000001110101",
        "00000" when "0000000000000000000000000000000000000000000000000000000001110110",
        "00000" when "0000000000000000000000000000000000000000000000000000000001110111",
        "00000" when "0000000000000000000000000000000000000000000000000000000001111000",
        "00000" when "0000000000000000000000000000000000000000000000000000000001111001",
        "00000" when "0000000000000000000000000000000000000000000000000000000001111010",
        "00000" when "0000000000000000000000000000000000000000000000000000000001111011",
        "00000" when "0000000000000000000000000000000000000000000000000000000001111100",
        "00000" when "0000000000000000000000000000000000000000000000000000000001111101",
        "00000" when "0000000000000000000000000000000000000000000000000000000001111110",
        "00000" when "0000000000000000000000000000000000000000000000000000000001111111",
end behavioral;
