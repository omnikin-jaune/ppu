---------------------------------------------------------------------------------------------
--
--	Pascal-Emmanuel Lachance | raesangur
--
--  github.com/omnikin-jaune/
--
---------------------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.ppu_package.all;

package sprite_package is 

constant SPRITE_COUNT     : integer := 64;
constant SPRITE_TEX_COUNT : integer := 64;

constant SPRT_SIZE : integer := (SPRITE_COUNT - 1);
constant SPRT_INDX : integer := 5;

type vector_sprt_pos is array (0 to SPRT_SIZE)      of std_logic_vector(POS_SIZE downto 0);
type vector_sprt_tex is array (0 to SPRT_SIZE)      of texture;
type sprite_textures is array (0 to (SPRITE_TEX_COUNT - 1))  of texture;

constant s_sprite_textures : sprite_textures := (
    0 => ("000000", "000000", "000000", "000000", "000000", "000000", "000000", "000000", "000000", "000000", "000000", "000000", "000000", "000000", "000000", "000000", 
          "000000", "000000", "000000", "000000", "000000", "000000", "000000", "000000", "000000", "000000", "000000", "000000", "000000", "000000", "000000", "000000", 
          "000000", "000000", "000000", "000000", "000000", "000000", "000000", "000000", "000000", "000000", "000000", "000000", "000000", "000000", "000000", "000000", 
          "000000", "000000", "000000", "000000", "000000", "000000", "000000", "000000", "000000", "000000", "000000", "000000", "000000", "000000", "000000", "000000", 
          "000000", "000000", "000000", "000000", "000000", "000000", "000000", "000000", "000000", "000000", "000000", "000000", "000000", "000000", "000000", "000000", 
          "000000", "000000", "000000", "000000", "000000", "000000", "000000", "000000", "000000", "000000", "000000", "000000", "000000", "000000", "000000", "000000", 
          "000000", "000000", "000000", "000000", "000000", "000000", "000000", "000000", "000000", "000000", "000000", "000000", "000000", "000000", "000000", "000000", 
          "000000", "000000", "000000", "000000", "000000", "000000", "000000", "000000", "000000", "000000", "000000", "000000", "000000", "000000", "000000", "000000", 
          "000000", "000000", "000000", "000000", "000000", "000000", "000000", "000000", "000000", "000000", "000000", "000000", "000000", "000000", "000000", "000000", 
          "000000", "000000", "000000", "000000", "000000", "000000", "000000", "000000", "000000", "000000", "000000", "000000", "000000", "000000", "000000", "000000", 
          "000000", "000000", "000000", "000000", "000000", "000000", "000000", "000000", "000000", "000000", "000000", "000000", "000000", "000000", "000000", "000000", 
          "000000", "000000", "000000", "000000", "000000", "000000", "000000", "000000", "000000", "000000", "000000", "000000", "000000", "000000", "000000", "000000", 
          "000000", "000000", "000000", "000000", "000000", "000000", "000000", "000000", "000000", "000000", "000000", "000000", "000000", "000000", "000000", "000000", 
          "000000", "000000", "000000", "000000", "000000", "000000", "000000", "000000", "000000", "000000", "000000", "000000", "000000", "000000", "000000", "000000", 
          "000000", "000000", "000000", "000000", "000000", "000000", "000000", "000000", "000000", "000000", "000000", "000000", "000000", "000000", "000000", "000000", 
          "000000", "000000", "000000", "000000", "000000", "000000", "000000", "000000", "000000", "000000", "000000", "000000", "000000", "000000", "000000", "000000"),

    1 => ("111111", "111111", "111111", "111111", "111111", "111111", "111111", "111111", "111111", "111111", "111111", "111111", "111111", "111111", "111111", "111111", 
          "111111", "111111", "111111", "111111", "111111", "111111", "111111", "111111", "111111", "111111", "111111", "111111", "111111", "111111", "111111", "111111", 
          "111111", "111111", "111111", "111111", "111111", "111111", "111111", "111111", "111111", "111111", "111111", "111111", "111111", "111111", "111111", "111111", 
          "111111", "111111", "111111", "111111", "111111", "111111", "111111", "111111", "111111", "111111", "111111", "111111", "111111", "111111", "111111", "111111", 
          "111111", "111111", "111111", "111111", "111111", "111111", "111111", "111111", "111111", "111111", "111111", "111111", "111111", "111111", "111111", "111111", 
          "111111", "111111", "111111", "111111", "111111", "111111", "111111", "111111", "111111", "111111", "111111", "111111", "111111", "111111", "111111", "111111", 
          "111111", "111111", "111111", "111111", "111111", "111111", "111111", "111111", "111111", "111111", "111111", "111111", "111111", "111111", "111111", "111111", 
          "111111", "111111", "111111", "111111", "111111", "111111", "111111", "111111", "111111", "111111", "111111", "111111", "111111", "111111", "111111", "111111", 
          "111111", "111111", "111111", "111111", "111111", "111111", "111111", "111111", "111111", "111111", "111111", "111111", "111111", "111111", "111111", "111111", 
          "111111", "111111", "111111", "111111", "111111", "111111", "111111", "111111", "111111", "111111", "111111", "111111", "111111", "111111", "111111", "111111", 
          "111111", "111111", "111111", "111111", "111111", "111111", "111111", "111111", "111111", "111111", "111111", "111111", "111111", "111111", "111111", "111111", 
          "111111", "111111", "111111", "111111", "111111", "111111", "111111", "111111", "111111", "111111", "111111", "111111", "111111", "111111", "111111", "111111", 
          "111111", "111111", "111111", "111111", "111111", "111111", "111111", "111111", "111111", "111111", "111111", "111111", "111111", "111111", "111111", "111111", 
          "111111", "111111", "111111", "111111", "111111", "111111", "111111", "111111", "111111", "111111", "111111", "111111", "111111", "111111", "111111", "111111", 
          "111111", "111111", "111111", "111111", "111111", "111111", "111111", "111111", "111111", "111111", "111111", "111111", "111111", "111111", "111111", "111111", 
          "111111", "111111", "111111", "111111", "111111", "111111", "111111", "111111", "111111", "111111", "111111", "111111", "111111", "111111", "111111", "111111"),
    others => (others => (others => '0')));


end package sprite_package;
